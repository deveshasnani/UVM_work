`include "uvm_macros.svh"
import uvm_pkg::*;


`define RAM_WIDTH  12
`define ADDR_SIZE  12


`include "tb_defs.sv"
`include "write_xtn.sv"
`include "short_xtn.sv"
