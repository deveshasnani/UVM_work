`include "top.sv"
// Code your design here
