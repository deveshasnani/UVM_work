`include "ram_test_pkg.sv"

module top;
  
  initial run_test("ram_odd_addr_test"); // try different test names here
endmodule