`include "uvm_macros.svh"
import uvm_pkg::*;


`define RAM_WIDTH  10
`define ADDR_SIZE  10


`include "tb_defs.sv"
`include "write_xtn.sv"
`include "read_xtn.sv"