// Code your design here
`include "top.sv"