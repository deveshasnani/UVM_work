`include "ram_test_pkg.sv"
module top;
  
  initial run_test("ram_random_test");
endmodule