`include "ram_pkg.sv"
module top;
  
  initial 
    run_test("ram_wr_test");
endmodule